/* Copyright 2023 (C) Peter McGoron
 * This file is a part of Upsilon, a free and open source software project.
 * For license terms, refer to the files in `doc/copying` in the Upsilon
 * source distribution.
 */
`define RAM_SHIM_NO_OP 0
`define RAM_SHIM_WRITE_LOC 1
`define RAM_SHIM_WRITE_LEN 2
`define RAM_SHIM_READ_PTR 3
`define RAM_SHIM_CMD_WID 8
