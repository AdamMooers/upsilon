module ram_fifo #(
	parameter DAT_WID = 24,
	parameter FIFO_DEPTH = 1500,
	parameter FIFO_DEPTH_WID = 11
) (
	input clk,
	input rst,

	input read_enable,
	input write_enable,

	input signed [DAT_WID-1:0] write_dat,
	output reg [FIFO_DEPTH_WID-1:0] fifo_size,
	output signed [DAT_WID-1:0] read_dat
);

ram_fifo_dual_port #(
	.DAT_WID(DAT_WID),
	.FIFO_DEPTH(FIFO_DEPTH),
	.FIFO_DEPTH_WID(FIFO_DEPTH_WID)
) m (
	.WCLK(clk),
	.RCLK(clk),
	.rst(rst),
	.read_enable(read_enable),
	.write_enable(write_enable),
	.write_dat(write_dat),
	.read_dat(read_dat)
);

always @ (posedge clk) begin
	if (rst) begin
		fifo_size <= 0;
	end else if (read_enable && !write_enable) begin
		fifo_size <= fifo_size - 1;
`ifdef VERILATOR
		if (fifo_size == 0) begin
			$error("fifo underflow");
		end
`endif
	end else if (write_enable && !read_enable) begin
		fifo_size <= fifo_size + 1;
`ifdef VERILATOR
		if (fifo_size == FIFO_DEPTH) begin
			$error("fifo overflow");
		end
`endif
	end
end

endmodule
